`define IDX(x,width) ((x)*(width)) +: (width)
`define IDX64(x) ((x)*(64)) +: 64
`define IDX8(x) ((x)*(8)) +: 8
`define rotate64(data,y) {data[63-(y):0],data[63:63-(y)+1]}

module odo_pre_mix(input [639:0] in,output [639:0] out);
  wire [63:0] total;
  assign total = 0 ^ in[63:0] ^ in[127:64] ^ in[191:128] ^ in[255:192] ^ in[319:256] ^ in[383:320] ^ in[447:384] ^ in[511:448] ^ in[575:512] ^ in[639:576];
  assign out[63:0] = in[63:0] ^ total ^ (total >> 32);
  assign out[127:64] = in[127:64] ^ total ^ (total >> 32);
  assign out[191:128] = in[191:128] ^ total ^ (total >> 32);
  assign out[255:192] = in[255:192] ^ total ^ (total >> 32);
  assign out[319:256] = in[319:256] ^ total ^ (total >> 32);
  assign out[383:320] = in[383:320] ^ total ^ (total >> 32);
  assign out[447:384] = in[447:384] ^ total ^ (total >> 32);
  assign out[511:448] = in[511:448] ^ total ^ (total >> 32);
  assign out[575:512] = in[575:512] ^ total ^ (total >> 32);
  assign out[639:576] = in[639:576] ^ total ^ (total >> 32);
endmodule


module odo_apply_sboxes(input [639:0] in, output [639:0] out);
  localparam SMALL_SBOX_WIDTH = 6;
  localparam LARGE_SBOX_WIDTH = 10;
  localparam SUM_SBOX_WIDTH = 16;
  
  localparam reg[63:0] MASK1 = (1 << SMALL_SBOX_WIDTH) - 1;
  localparam reg[63:0] MASK2 = (1 << LARGE_SBOX_WIDTH) - 1;
  
  
  localparam STATE_SIZE = 10;
  wire [15:0] next[9:0][3:0];
  
  localparam logic [8 * 64 - 1:0] sbox1[0:39] = '{512'h3C2D3F0A1A210E033E06221C392C2B270F162A29341B202F383D2E04050D3314353B3A1801191E322337131726240C0011151F10311D28300708253602120B09,512'h020F142D1C3E030A2739302A232429051116181219062C361713350815321E3F3C21000B343A3B1D2E371A26042B220E20381F0C281B093D0D0131100725332F,512'h3716272D0C11391F1A323305252F311C3E2C1310342E303521023F29031D3D150A360100061817282612243B1B090D380F193A0E3C1E04140B2208232A20072B,512'h3B1F332C282609203C19353E042723113A24130806032A1C071E1B0E32223F15300C381A18363D0D0B2E31001D21372F390F1714012516022B12340A10052D29,512'h0E213203373933382023020A08002B3611101407222F0F1E17160526303F3D012A3B2412311F1929272818350D2E3C3E060C2C090434131D0B3A251A1C1B2D15,512'h2A352B360F3F1708110034281A30371514291F2D2520010921022F0E1633123927193B243E1D063C1E03182C323A0A0C1B22230B101C3D382E05040D07261331,512'h3F200D261B3E2D3C001F280E3003171D331824320201052C141A2E273711210F04293D090B25133931342B380C1C222F3B072A19160815103A35231E060A1236,512'h101629041A3237173A1E190521002A0130023615223339240E0A2E2025110F0826063F2C142F183C3B12340C0B2D1C2707133E381D1B2B35033D091F0D312328,512'h060B112207163210010F2B2638281D1F3C1C0318133E191220232C092F0A151B3D2E252924390D21173A3134053F2D2A353702000C083B04271A330E3614301E,512'h1525052239230136373427320D20180E28190B2A1D3F042E3E073B3C382B351A061F09311213023D0A170800261C291E161B30112D100C0F2103332C2F14243A,512'h1131260E201328010D22231C031402182F1D17293B1007122E0515323C3934082B3506303837363F27211F1A0F043A3D2D1624333E19090B1B002A0C0A1E2C25,512'h2227022C3411231A2D3D392B14170E13253F20312621060A0D19240C10163515322F0912071D1C03011F3630332808373A0F3C2A1B3B2E001804380B1E3E2905,512'h3C2C3E27382E02191D0F353A3304281637312A0005361F1A1C153B010A32233003102F34070E1E1B183D2921111739090D122420133F0B2D2B0608220C251426,512'h2032212B2C091E06383E270836121B3C101F052F0E0C340D133914223035242E071A0B312D3B1D2901040F003733181C3D3F261123020A2A281625153A191703,512'h33362B2D311D0A2307132A0917242200111E342120123906143E0B08283C37040F3D1926181C102E3B1A29301F0E1B15032C32053F2F0225160D3801273A350C,512'h32010214380330251835001E293B130D15310B050F27330E2A282239261923110C1636123E200804372F3C091021342B241B1A071F3A3F0A063D1D2C172E2D1C,512'h3E0F1D2C382831142B1A0C123D0617091B392418163F3C2F340D2730291C19222625352311370B3308323A2E2D36040321021305073B011F1E0A150E20002A10,512'h340510171D183015011C020B2108243329231F3A2D2A1A2B1232203F04392F370E1E0309350F271B313C0C160007133E112638222C363B0D193D2514282E0A06,512'h2B26090C2A3A162D292E3E0F1B3C212012112F17181E3B0A01032315241A1F193713003305311D283902361C0B0E38223035320D270806143410073D3F25042C,512'h0A0036340513063F18333B171A2026310824270B3E351F2E2F37071415321103042D0D3A250128290E0F161D021C1E192223392A09212B12103D2C300C3C381B,512'h161B2B252E113C27171E3D100204232F1238242009362914083B1D0013070E190B28063E18322A1F35153A0C300D3431053922332C26031A1C213F2D010A370F,512'h2B0F020B041D090528062F08181C1B2E0A1A3820321437133C3036073A1F221E192133352A3F29170E251623003401113B2C3E0C0D102D31242603151227393D,512'h043C3B2530262E201F103735321614191C292F0A0D09281303341B18051A0F33063F112B231D272D390815123E222A000B1E360E0C3124380121172C02073A3D,512'h170A0429241D300B0E083D15112F3518223B072501061A2E191302380D3A3C05340F3714231B0939122716200003282A3E322B261C3F2D2C1F102133361E0C31,512'h022C090D2B393408191D063818353E2621281632041431002E2427010F300C1A1E22053D2A0A3F172512362011101F2F333C1B072D15133B23370B29033A1C0E,512'h1F3F033819053417210F333D223E150A02391832090E23112B1E0037160C072F1B2E2520142635013C0B241C06120828043A1D132910302C271A0D312A363B2D,512'h03061211040C25373E22021F3433392C362F1810143B1D1E010729161C0A172B15133C0F383F2A211B2423080D192E3A003505262D323028273D200B09311A0E,512'h230B22313B380A302A0E1F1316141B32090F2F07051106243D100D1E1A36041235372603252B291D02083A2E17192D1828273F2C0C1C15000121203C393E3334,512'h1F052432193E28271D3D0709303F2B1017313A3C340A251A0E200F2D1B233815010326111E29060D35333B2E1C0416132A2C0C021439360B372F122208001821,512'h0B0E0231043E141C272F12010D2B180F221E30103421332015051D253C1A0A3A35261B280C3707133608292E090600032C3D3F241123381F16192D32172A3B39,512'h0F012C3A2F280818133534220D1A3B2A1D14001E252E120A1F26382B37031921070B321B0E293C3031041C3909360520061023173F2D27153E243D160C021133,512'h0229082107351F033E260A3113002422341204052815103C1401272D11230F1D1C2A393F321B172C0E0D1E1A160B2E062B3A3633253D0930192F203B18370C38,512'h051D2D3A02220A2E131916030B271B091C3926230C2A3C38363407313B3F0D3D17182F1A0425291F332012061015212B112430322C0837140E3E0128351E000F,512'h203D020F38072B281F120325163A0B1C1A372E19303C0C133915230431052F34002618213F113332171B060D09360E243B291427351E3E1D102D2A0A2C220801,512'h04302A0D0222062D2100201D083B310B1A05241E281517331338193D3F2C0E2E390125100C18361F35343E1B120A2F071C030923112632370F3A14162B293C27,512'h0B030732133C2939001D283534023B052B37313D091B21382A193F2E201A360F270D1115173A231C3E302514082D0406180E24162F0C0A221E0110122C1F2633,512'h271817191D30321408212A3931162D2203342B3C3604000B2E28070601151A11090F2502203B3D1C35233F1E123A0A0D263E0C38132937332F0E10241B1F052C,512'h2215300110022D2016333E231D3C313B180E343913362B083F270C25050A04061B113D38121C2F19031A3A1421170926002C291F1E2835070F0B32372E0D242A,512'h1D260D0813170936242D2E0E061504300110023B0F2B190C1F23222914123E320533181B3403000A3F3A281E0B351A3D2C2731252F382107393C37111C2A2016,512'h0617143F372E05040A1D233C070E090B13280F0C342410191C292B2F1E001B1511303A3839350D3201121626223E3D3B2A25082D021F20212C1833271A313603};
  localparam logic [16 * 1024 - 1:0] sbox2[0:9] = '{16384'h00040191014A024102B102BF013302A90147004701F8024C00260178022201F202D701E201740295008C034701FA019403A8024A01230358003B004E0312019603D001A700D400D2025A005002CB028601B4012F035503FF0251015B01690395027E007A0392037703E5036100AD0027015001810053009F033801E7025D02A2025F03E901CE000F01FC00010253002B001A026F03A7018F02D200A20352037F03AB0151026E01B800EE013B02C201EE0278026D0382010E022B02EB007602D8028C02A7003603DB03CD013502B70052020603F301A3019E027703E700EB0089037A03FC02320035015903050385032200AC02C7014D0331033903F401F4014E00A803C5033A01ED0254029700A9003C02790144001902FF03DA020202E3030000A5005D0289006403D902920018000A01AF028B01E900F1001D006501650242009B01290183002A0038011E003F01F602B603EF01B003C1009200DA01E8005901BE011B015200E4022A039F01A60266031701320281034F02AC03900085021E029D013603A503BE000E000902DA0011034B035600B3000D03B902190243029C023B025B01C60272009303F0019502690200011300A101D20043032F005E0197035E030200730369004502E10209012B006A020401EF01D801E503500258034E007203C3008A0367035D03AF019A02A30217015D02F6019801F1027C01A4002002610055008B034C00E30090012101D10125010600710237019303DE0006030C006B0057037203E001C100C102AD00DC0008018C020B022103BD03DC024701DD027102D500AF02B80255006E032900D0010800D8019202AB013003B40216006002F2012C01C903340112009802DB029801E3031F00D100C203FB00BE01D900B103430330013F02EF002F0393008F0134025603F10013018A0137002C017E0139026C02F502E2021D003D00F8008401840205034002E60324007C0267039E03B20079007B03DD03C003650002031901FB03C9033C027D039801EC01AE01BB003103FA02DE015802F3017A02DC038100A4011F00A300DD0366034203E602F9030801B7007D03B801DE02B3021801D6037E00C5034D02EA0235011000C00287013A03CA02A5032B03FE000502880321021A02600142035702930030027403090229032D006C022402BA018D023F025001E1009C0154013D00560388038A0170021400620083039602AA004602D600A6004D02E703EA00B6017F022D021500ED022702D3029F026400BB024400780201006103D301FF0370013E03A401DB01C8006701F003AE01E0008D020A01CB0211030E0087012D00EA038B0171010F03140153018200DE03B0022C033500FD0228029900C3003E011C0116001E023302F100B70383010301A9008000E8026202FB0104031E016C01D001AA02CA00F3020C00F402B501DF03490375014C00FA0012009E00E2007F031300E5017B033F0245033D00150208018B037402D9002401DC03D10310010B00FC03C2038D0160017C030D0016035C01D7039B037303D80384010A039D01C50146031D03E801B100BA016B01A202C303FD024D02BE027A01AB00D502C601C300FF0145030F02DD03A20231024B00AE008200400115004202B9008100F9003702F80179029102A80304001F00E0037800EF036002CE00AB00E101BD02A6024E019C010C008E000B036F027F031B0362035301C4022602B402AF01660270025701CA02030105028D031A00F6000702CF02EE00B003AA008803D60187026B023C02FC00C70186020D037900CB02E400C602B2034503C8006F0380002D014F036803B302C80265024803E100F201A1019D0094004B0315025901CD0054029E0364005B01630017017601FE018801DA01B302BC0234036302B002A0015501C2016701B5038C01CF034403C4024F0101033200DB003402BD00DF0138018E03A90225019F001000BF03D500B5014103E20391016A037601A5028F024902D401D403F6002E01BC033B02EC031603F803BB033E00CF03CC01750095020F0268027502F70048016E03D701A0010D011D02ED028201E600D7038E023A007501090189007401A80033039C023901620120015600E6028400BD0102002100A7033301EB02C003A302E5034A01C703B70131035100C8015C03F2032C030701BA036D0023017D02FA00C40246018503F5003A00F0007E009903EB026301640086011901F5015F0290032000960311032500D90190016D03CE037C027B00B8025E02D103B5015701D503030025016F02E00000024001400127037100D6021C009A00FE025202120122039A001B011703F70143016100B901CC00580100012800E903A0023D00FB01FD001C02CD0091032303180210020702BB03B1011A0077005A020E028301BF00CD03BA018000EC015A014902E803CF03A6025C03A102DF028E02F402AE00A001180049014B029B001401E4036E00E702FD028502E9009D01F9039400F501EA0111030B033600CA029402C401990348006D03CB03D2030A00D3036A01B6029A00B20044034103E403280003015E023603BC023E0097037D00F7019B032601260397022300CE01730068022E005C004102F0012E02A40051007003DF03E301AC01AD02C500BC01F7004A005F03EC0148003902FE037B006600B4030100320399013C0172000C03D400AA028A0230027302C10386029603BF010703370213021B03ED004F0238027603C703AC03C60029006303270220032E03F900C9035B0387022F0022035901B2036B017701D3031C02800114036C026A035F02D003B602C902CC01B900CC012A034602A10028032A0069035A038F0306035401C001240168021F004C01F303AD03EE0389,16384'h001302A902C902DB025603CA02EA03AA0036017803A9017001A500F6026801010065037D029002E302CE02D3028F02E1005503E900E1004B00FC03E2010201CA02F6023D039803C2002C039C011A0298012A008C027000FF008701D703600356020F03E002FF035200F70035019800DB02B300DE01FC031001E80306039901D000AA010703000377016903B5034B0348007703B800FA03B003FC026F012D03E503EF018103CB01A001E6019F01C20081009A01BF01280097015702A003F100540201019E0094029D03B301D300B0021B0005012B0243019602230251037C03AF0183036E008F003B0009015A01C0000001D803BE03A500E601720343005C02C100E0031B00D6020C015303740112030E015103FD018201ED02A1030A03DF013901A3031301AC01AF02330190027C0056028101F702F1036D023C019B016802CB00580369031A015C0173002502DE0370021700700323024503A2015500EE026002B5011003BD03BC000F0390032E031200280350018600C90331032A0273006E0003026D0048012400B1024101420293031F020001D601AB007F00AD017B02D2002E0031015902C6028A027500BB032F0368017500B8008A00C300A103380045026C00D0022501FF0068001C037903F5038200FB0160014C01D20396035C015D006F020D01F102C5017C021300D300990309011E01440105020703A802380002032D025C02A401650286002B03C103920162029E009C02500292031E032402CA0206006003910333039A01BA01790364021E0287025702AC01F300610088026E006C030202D8026601CD01A80029006A02D1039503F3037500CF025B0325033D018700D7001700760113034001A203C600BD019A00780135034A00B9020A0176002A0239028C00DA000D0262034F0376007B02ED0214007500D9021100C8038D03C402C002BA03EC01BB025E010E0026022703F20278031C03BF00A601AA0285039401E30276030800340171026A001E00E903DC01B3031100A701C7035E0341011600A4023100B701B402480191035A016602FE02CC005103ED01E2015E003902EE01A90321010B0103007C00DF0147015F00F4018C004A0082022F009503F9027A02FD027102E9024C02EC037800B501460279023F01C502DD01DE01EE0314021F00930205008B0161022901D50299034C0336009D02020261012000F1014F016E01C602F2004D029703D001E701190092026902D502EB00D10184008E024F036C00AB014B02E803B7027202EF017702E20064014100BA0106002400F200BC02B602C301F6021601B000A50156018D0083020303C70282014A03DA00E2032B03E702BE0235039E031500C5037300CB00FD013F01C90366008602260118013300F902F40264017F00DD038102E6031702B0033A00C7001000CA02440137038600B4030C03A4009F005A02D000C001EB035401D102F8003F0346038C0265038000C1029B02550210013C02D4038301B7035D010C024A01C401A102AA03BB00D203010041016B0236022200C6028802D6033F01CF01220038011D01E5019902AF01FB00C2026B02FA003C029603CD0030000B03B10138032703190132012E023B016403FF03B203D6011C019301EF03D80259034E011501C8028D033E03BA00470384035F00EF0316008001DC004201D4001D032203E102FC012902F301EA01E4010900D803DB02670008007A02F903C0033B033901F40185003A02D703E30234018A0014035100A2038B02950228021D02A5005B001201CC02F700BF033C02B2007103AE007D001601F9035503D903F000E70209021A021C03FE0040013B01BE007403050247011B022C0304012F001100B202B702C8002D0043005F03DE03B602DC02A202BF019C017E0023002101450294000101DF008402E4001A01F502B8022B009801BC022D00670050037103C8011402080318001B03CC012C018F025200CD027F00AC01DD03F601A402BD03610019025D02B103EA036A02B4002003D1023A01E90224024200F500F801EC0326002F01AD01D903CE005D00A801A600E300630180030D01CB01880397032900FE03DD028E009B010D00A3016C01FD017A00ED0126037A00660328035B0123030B03D40096025A0307038A0393010A0232021801080143012100D50027037E01F200EB004900BE00F30365028401E002E5018B00620085001F025F009E02E7013102D901B500EA020B03E4021501AE0388019D003D017D013402B901DB02AD0283023E039D034903EB000E00EC035302BC0344021902A30230008D03AC026302C2000A01C30195000C006B036B029C011F03C303570007007201270117038F03A003C5005201300192016F00B600F001DA027403AD030F004E016D003201BD01CE03D503C90363001802A70033007900AF01FA0289001501B2032C00CC03A600D4013A028B01250037029F003E00220362023700AE03D3024002AB016301F00335027B027701110069013602C40148022A0387033701B6005E00A903CF016703FA016A00E8037F020E0320010000890280014903A302DF03E600C40367034501580246007E0140024D02120194015402C7033201B8010F02A802AE03B4033002BB03720152013D01B903D203340220019701F803B90004000603F7009103F8029103D7034700B300A00073018E03AB01E10044018900E5014E020400E4036F025802F501FE034D02FB03A7004F0221004C013E02DA0090027D014D025301500057035901B1027E039F03A103FB024B005902E0004602A6030303580053025402F001A7024E034200CE006D038E015B02490174031D01C1022E02CD029A02CF03E803F40389039B03EE0104038500DC037B,16384'h006600450192019B02DD01B103F002C30220016501550252010800CA00F60310004203400017032302ED02BB012F008703E7027F009A010D031801240312028702C0016B012303A602AA0083020401CF01A90359005A019C004C0036006702530135020203FE01A101B803AF03A1000A00AC036B03E1005D03B603CE02AB00E9013E035E01E503C7014601FD0363031F00C70217021301360221028C03D901A202B50365024B0182024501450160002102E700110004019002FB00DF01180244033A00C1002D01830327029E02A4003B027A0360017C03BE029502AE01EC00DE037D000702A20211004F016C0288032503BC03B2009901670030038802620330011A000D00030158012B03B900400041018A037F00F900E2034E00D500C60396002B01340358008F022B00A2020702E8002F0001032201D902D402CE020F02CD0335033C028A00BA02B30088003A016F0140036F005000C003DD037301260035012D00AB00E7014B02E2024D013C0053022D021C008101BB02B802DC031301DC02C803F9034500B0019E021D01C20255009403D803EE025E00D6018F02EE021202FC038B01F6013703DB03A3001E0387022C019703F20339025D00B90065016D0385000C01D80303019A00E1034902B9017D026503B0030C0082012000A6005F010E039401FF011101C003C9015A006B01130070033801D3036C037403DE01AA0080024C03BA00B7039E02D8015C0060029B00EE0379023E021B033F01B7030D022E00560264038601270199036402F302BE03BB024300FE00CF000900F703D00191010A006103F4000F001500E4026D005B033303AC03C60368002502FA01CB02250095029F032C026A0059013302FE0144027300BF018C0397020602BF025902F9003702D0018000980141025B03A2017703CD023701B901F0011C01B4015600AF036903E801EA007B035503E603AE03B402C5033D01320376008900B602B1034D00FF037C001B02CF03D7015D022A017A013F01EE023201BF01E2028D008B009B0301035001A7004B0052013D02500239021E01BA011D01380149038E0246035F0294008E01420271021F022603D2039103B30251037800F3007602280343004A011E0006019303E5001A00BB0296009702DE018401C701D70278025A024F0308026E003C001901C3009103E0019D027500F800D401E002230254025603200332005400E0002A00EB03AA01E1032D02E3006D02CA00E60196003D0331031A00280281011201CA032E016E009C0031010C0277001F005C00EF0361012C008C01A5000500F103FB00A80304002601AF0139029D00D700DC01B5039C039F03D601E4017501BD01FB0305022202D5015102B20382034F03F8031C01700150028402B0034701FC00140115037003D5017300AD039B02A101D10276001D010703ED0297019501A80178023803AB008A00A000B300F5026C0293006903DF007803EC02CC0356032A01C80103021903F3005701EB00A900B400CD03F5013100960392024E031B01300267005E002E0048022902E100AE03A4011602D903B80342017B0121028E023102E00214026B01F8002C0352037A018B03C103A5038103A8032402AD00B8029A02100274037E023502A500ED00E301B302B60234017201AE03660162035701C60198017403370068009F032B01ED01E600C201DF03A7038003950104023C00D2031E00FC036A000B02A803150046007700100148002000D001A602F0010002EF027203DC006A012E00A402980171004900B20283039003840166020D038D02A0018801E303FA03E203E401690269001C00FA015201C901CD0309013B0346001302DB02FD0216023B006E031101F2035D034C016103F702EB005101FE035A025702E4006301C50117022401A0002903B5009201020285028F0336022F011F034403E303B701F100750314014F035403C80247033E02F203CC032902F100F2013A00C300D901CE00EC0110037B009E0002032102DA03BF027C007E0208007D027D00270128026600DB02E502580085014C02A301D20187009D0292039801AB03F602C103CB015902C7016802CB03000201002203EB02BA012200BE015E031603DA02E6002302A900B50236006F012A034A036E0249020C0119018D02F50209015300FB014A01B0008D03D3010F0279034B024001010106007C0114030B01B601D601E7020A026F02DF02AF01F3023D02FF007300DD00B103CA03FD00A1007A035C037700EA0164025F00CC0176018502F70362018900D8037201F903CF038A00720389031903C4027002330334035B01B200C80163025C02420280020E039A01F501F7036D01D0028B0086010B00CB01D40071015B018E01DE032F01DD01C101BE017E00C5004E03F1002403EF02A6014E023A000800C40268009302990291003800AA036700330375031702F8024801CC00F0011B00BC006C003F03B10227038F03C0028202F600D102D302050034037103D40383024100C9000E02EC014301DA015F038C01A401C401E900A7004702B70012007400430157005500DA009000790348027B03D1003902BC02D700E8023000CE032603A902D201810261027E023F030700BD0290032803060062004D00F4020301AD015403C30147030A02A702C402C90016030F0351003E03E90186034100D303AD0032039D031D03BD012902E9007F0194020B02D1033B0125021502C203EA028601EF016A0044017900840058019F0302035302EA0200026301E80105000000A302AC0018021801BC00E503FF01F4026001FA02BD03C201AC01DB02C603A000FD03C502D60399014D024A006403FC02B4039300A5021A017F0289030E01D501A3010902F4029C,16384'h033501FE027000DA0329012101E200730387004F01EC026B0233034E012F033002C4008001AC0025037E027700BC016B02FB01B603460326033D00F6017700D402E90378014B000401DE00D70358015C002902B7038A0149020C02F1033A01E40251012D0371017402F3018E0155038D0286021302090009004703E000AC0065018F015E026A01C9024D03AF00CC01590287038203A80385013501C5037B007A00F00267019201E702A4036B00D0032C010E005A016F0176024C00E203A90237031D03BB03C5034F03DF018800B4012900BA017E03D6034001BF00CE0052032A00A3001C00B703A602B503D5019A03B5011D02AF005C0144012800060216007602C20136020502FF035402A7011C00EA01A7033B0112000201ED035D015A02DC00F702D10003005300950070001E02F402A20057026903B601CB019C03EF017501F900CF0199029D003B03F30039006C02FE02F603EE00DC00D200AB00D5009600B10141028B03DB03C1011501DF01AF037701F603D10161023D00D9031F001702600289009C02A8012C029900A801200381006F001A0242018D006703D303DD021C03FF021B031602E000E502B1030C02C501A3023602E501E500FC031A002A0215006A0271029203660322011401EB00C20344018602C8003F00B80365035C02B303AE00C102D903A103CC035A01BB003300B6014D01F4020A022601EF01780042038E0173004D0353022F023F013C016E01A101A601FD00F301FC019301C102AA03DE028E014F000B012A027B00F2032E02B20098017201EE010C037400BD027402BD00900093035F036203940030013300E9029701E6012601FA002C039F039A01DD02E6023C028D01950171027C00C9003A024400A4017C037302210181002E009B008A011100A702FA0259016003BF0245024B0132006E019700D3001B0075008E011902410185027F03E80005021A01D200630069004B007F010400FA035B017B004E0285017D033602730243008D01CC02960170027902180194014600790338030701CF03EA02AD018B02CD0048003402DF016C03FD0084024E034700BE00C5014C017901F8039B03FA029C03250072002F008B013702E30145021E004101F703D8014E02780058011F00E80229032800EE0312031E0142011301C3019F01D000B902EC0261031B012302DB009A039502EA0256037200DE00F90180013E005403BA0284021403C7002D03C602D7039002BA032D03A7021001BC03B402F2005900CA00AA013F031703FB02A5030603D20086023503BC0211007B015B03CD030803D4002003F20026038902EE01DC006602AE013900FB0165033C02B002A001670038034B0014031C028A02AB006002E40268025C01A900F4030501EA00A600D603E203C801D5009E006402CA02D2015F01D8015601660230020E0290015203130157003201E9005B028802FC01AB00CD015000C301FB02030350034D0337026D02BF030F0240025B015302980281033E020701A80263021702D601A2021F02A600EB0282027A038400C4010F02FD03B00044039E010B03C002DA0383025F035E03DC00ED03A00396022A0013025A00990352029B006102A3005D01F203A300E403F10081018C012E01C8004502060399022401890319033F02BB01A000AE007D0021019E026502040083001901B003C2027D03EB024900B2029402530012029100DD0272026203E501B4023A039702EF0049001503D003F501C4016903D7010603BE03F90304004003BD026E020B0348009F018A03B1013800A002A103E9028302BC0140038602C303C902E8034103ED022202380388023401B90028039201F30164036700FE00780368016A008700EF01BA02000295021D01180122033400F10125023E029F00CB030E019603CB00DF014803F601D903DA01D30332004301D1025000E1009703A5020D0247010D01AE01FF02E70001012700370184037003B702C903210101004C0085022C00710225010800B001870252000E00DB0011029A03EC03910088009D03E100FD019801E101B7003D00890355012B000C006803B9027501BD026C03AD01A4031400C703450050001F01F1036E038F02BE02CB024F00240110034A005F007703D900A5017F00510228028C030300A90191003E02CC017A019D0300035700A101E30007021902C600C80351011B03AB00000276030103100212027E031102C1036A038C02B9022B0364039C00BF03A401470302030A03E600E702DE01C203E4011703FE01B5000F01D6037901E803E3022002A9032F037A03590154020F0201015D0363013402800130013D029302F0006D02B6014A031802E2028F005E038B00E3007E016303A203F401CD039D02C70361031500A20105016202ED0343008F0257013B00550223002303F801F0025500F501DB032B00C001D401F5034200BB02B402F502CE019B009400360258000D02B80046008C02C0025D03B8034C02F901AD024600B503AA030901C0004A011600B303CE00740107015803980266013A0232016D002203FC00E00231008203AC0182010A0320023902080183006201DA03CA037D0254001003F0032703E7010302D501B1022E011E01A502F80091000A013102DD03C402D80151003C029E001603760360037C034903240380033103330375006B00F8001D0056036C00D8001800E603C30202002B02E1030B009203CF016801B8003501CE0356037F00AD0227000801C7012402CF03B30143026400270109024800D101BE01D702EB00EC01AA01C603B202F702AC026F00FF024A022D036F033900AF01B301B2032303F7030D011A036D025E0190039301CA01E000C6023B010002D402D302D0007C036900310102,16384'h004702D700D3038C022D0372034C033D030C024C03470249014E02440166027E02BE01320230016100CA0231031503A500AD030F00D7006A01FF0064030103570246004A00CC0107006F012701FB0362000401D601C70211000F03C103F101AD00C90272015402DC001601C3031902DF021300AA03BD039302DB00EC00580153002800C200650247010E006603EE0100004800AE025C033A02920371028C005E02A403E2036F00F200C50332036303F7011102DA00BF00B9030803C500BE0136014F0221010A01ED0388010901B101A0024A0157028B003D032F002B017D01C40134027503FB03480337028D00E9009800D802F603200138032B00A1027C03AF003A0288020A003C0181017B03030199020D006803A3034001AF039E01E701C601CF026B02740309026A015B03BA0359034B018A025B03B403F401AE021702F503F9035C03540305026D01100141000A01F1038102D8037C00CE004F00C30080032403CE0148027D02E903EC028F02050019026102B1011C0234029A02F801D000A00210014D02D50059002103FD03AD0365012E011201F602840334033003C0032A004C00960008030403DB03A0014301B300AF03830240023D0018031101E2024502FE003B0346029C03870214002703ED00E4026F011D012602F702FF01B701CD031B03E0038A03D6008C0265038D00D1029001CA0085024802B90239018D004203FF034A035E0218006C023E0034018E028A017F012A02C403B5014701D8011401AB02A6035A00B2037A017C039F01DE006E03FC02D000870123027301EE00B7007F03FE02AD03C2009A01820145016703B801AA024E01C1014902A300A602AE00EB0131010D011E00E7009D029700A5022601020256002203CD03F003AA01A701DB0188031E036C01DA008E03820294023B00CF00F402F2004D00D400E200090128019002C200FE013B03640049031F025E032300C4001300150093012C036B00DE014A019A01D20017017801D70390027603170328015A01FA020C02AC03E9019B031A0037023A0144029102D90129013C02CB00F302AB02F9010101F902FD015F0030031C01650258002901A6020E0089000D028902B501A200430263007A00FF03A4011A014C01B902CD037E008F02F1013A021B025702B301F50267022C03DE01B402B6009001E8039803C9033E039C00A8005F01DD02BD0227028001AC03D1006901680158009C01890336007D007C0014031D0045005203BF0314020B005401460026004002BC02D100DF024100B00243007801740216011300ED03D802BA03EB036601FC01930175024202D602A102E6036A03890202018403EF001C02150036021C0120017701CB02F002C7018501F30338006D0024002A03B2026C0135001D029D002302600232017603DF011700790039039702EF0055013F03B10250027B001B03B60350030D039502FB02D200B102FA03350306028501CC022500830327003101BB03C602A800D602E20386034100EF03B003D901620061016903E400380187018B000B00A400F00352003200A200E10091012B00D0038F03A200B6035500FC025F01A1038B02EA0344022E015100C7005A0086012D01BD039900DC03DA011603180041030B02CA015E0001026903BC01A803B9021F02510160033102D3002003C8005B03B7007202350307011501B802000361035100B303E800C0016F02CC02640300036702090392000E021A007B01F802BF033900E800920171016302820005039100E3012401060198012F03A700EA022A00CB037002E002F40173026601E402AF015501E30033019E023601A3019400DB017901F2015D0046037B003E02C501C203D401EB021D028100500296005C02D40010008B0002016E00A901CE030E032E02EE0122007702B4001E01BA016A00F7019500E5029E03C7033C02E302FC033B02E5025A02C30356025D0074019D01800259006700BB02B8011B039D01B6011803A9007102790073009F0172002C032D03CA02A0012500A7005101BC027A01FE00D501EF00DD02E8029500B803BE03DD019700F6038000C1005302A50322020601BE031200AC01D502CF02C9024F009900E0039B0349037F022001370088029903F3026E03AB019C0035009500F50378037D000C00BC026203E6008202B002040108010C00C800A300FB022401D3001A01A500B503AC00F8013003D703450076011900B4007501DC032501B203D0037403A1016C009401C50254025502A902C80000020F0152023F0170012100F101F003F602DD002D03A8032901910007013E028E021901BF01D902A7030A03C3034E018301F4010301A9021E002F010F03E102F3009703CF01040003022203F202AA022B003F02860233016D028301B5024B017E0310005D0044008101FD009E01E0013D026800AB034F036E0006035B03CB00620203027701E503D2016B011F002E0394020703770270033301E103D301C00156009B022803EA00FA0139027F005701EC01920384020103160278032102EC006B038E034D00BA020800CD03BB035D03E5018F00C6024D02E40369039A002500F9019603C401DF02EB03E70379035F00FD02C6018C03A6029802ED0105001F03130343029F023802C0030200EE037302DE02930056004E0063028702BB03F503FA035802520140022302C10011007003DC01E60353013303F80164032C03960060010B0375007E01A40342017A03760253008400BD03AE02E7033F036800D901D400D2021203CC029B03B300DA019F02370326014B0150015901F7008A0012015C01B002B70360022F01E903E302A203D5008D02710385018601C900E601D1014202B2036D01EA023C004B022902CE01C802E1,16384'h005503520004033603FE02FF00C9011701C5019703B3005B0000031200A1013F009D003900DB038800340129021201BC003F02AF0081026E01B702B5008C02A903FF024A007E023303CE017200EB0191014703D50230030F017302FB032A02520035021B03A502800185035C0224018F011902DD039E03A8002D00C202A7013903DE012702BA011203AA01A8014C0097005300E201B8016F0295010800C10064010002B902C501260257038C030603470346014902C0020D00EF029602F703A2036F014001EB024F00C401E5015F015200C8017A035001D30138018702FA0136029000E100C602320171034E02DF019203C500520254011C0181018A01EF00FB01E00365037C028B02A002FC0303012002040248033D01AC020203F8032D03F6002F017F01F7032201F100A5016A021C0387015B037702220276030B01C6004E00D3009A01A90269010602EB025B01F302590376021501FA0305034F004901CF00F402AE034400FE03B7039301D101D903D40372022D01220008010C0162003D022A03EC00FD028A00B6039F01F901B202C402620325002903C3006B0239012D006001F003BF01FF034803B80194030C006C01A7004B0373009003BD0105001102830301015401A501E90340018E027F01630357002A03C201DC0379017C00CA004C0088019E021A02B1026A032400F3033E039102DC028D01CC033202E0016B00A30072031B01EC02E2039200E8038B03170319030A00BA03BE03C90333000B0397008F03AE010900B400820094003203C6022B03F203D600AE000203C402E701DA018B02A800BC013A01A203FD010100300165000A010A039903940238022501F6011F03D1022102E402FD0209019802AD0263015D0047019303B600D1007101E300CB01160042032C01C701DD02910211037D01BA00BD01C4035B015C034D01B403A1001F029302C10123016D02F8004800590045015600ED0264012801AE03BA036C035F03CC025600EE00E502660155031503CD0043005C01D20098013001C8010203F100E6020E026D03B501C901D0026C012C0118002100B50115017B00F503A00027021E0174011A01B501CA025C01F2013C015900E302B400FC004A0251008E031800A4032102A401DF029902B001A003040300019C026F037E01C303F300DC014202BB023B023C0038002303FA03F500C003430383036D022803D700DE003E029C020B027C030903E402C600A703B10345017E02C7022303690335013D036602F9037B01B30014039D031C028C01E2027902860307009902BF02EA00A9020C028502C30292000D012B02DA039B0153008A00A601D4019503E7002E020102C202D203ED03F402260012009E03F0002B0062024502D90288000603300075020003B0038103C8011D0084019F00DF00F103D3007B025002F302BE010B021000E700F901F8035803B203E30243007D032000780271025502F403750024001001D800CD00B901E80058027503EA0124002C013702D002270151009B037A01F4036303C7021700C302C901D603600208038F008D010E02970066029A005F0107009C03F70287017D001300E001C10184026803AD036403A3019A02F0039C01FD038A0168013203D9025A00090085036B011B00D503BC0359027D03E00362023100CC02EF01C2020A008003DD0196004F02B801FC00F80390011300D603A70199024B023500B001BB00B303E902610141020503610057001903FC0207033C0033035E007F001C00F2035D01AA0281020303DA036800D2026703BB026502E60310038203C1021903260384028202D601830234010F034A031303EF02ED022F025301BF00D700650308020F038600AC028E00C500770374024701500091025F03AC0258011E01B6035502420050037F0157007C01A1003102DB02CC01EE023D03B903CB01B1031F00A003DF0161024C0380006F00950103021300FF0339029E02E101860327019002E8013102EC006E02A601F503FB02B601E70370012E038D02290114034C01CD003B00AA014501660007008600E902F5005100B80067015E00870342004400A20398038503D202AB00760272022E0028018900680061028900B2000F00BF007002D1029F0040005603A9006901770083019D02F103A6008B02740284030D00A803C0003A0329035600C703DB024900E40294012F03E103AB039A00AF022C03E800CE03D002A500D901AD023702EE000C0180026B015A02D400D002A201AF0017030203CF032B0104021F00960164014F02A1027E005E03F9013E029B02AA039501CE0073031E036E0214016001B003A401100018005A02440005033A027002E50092001A02E300DD023A031A021D02E9001B004D002201AB013502D703AF02D8032300F7001602DE0167001E00BE016C03E503E201A3014E01E6007900FA02D500F0012A02CB0241012501A401E101780020037101C0007A02CA005D034900D80025013B038E007402AC00CF016901790273033100F6033701A6012102A30170019B0378035401D7031D01FB0041000E03EE02CE02B202B70054006D006A029D02F60341014600AB011101820353034B00D4002603DC032F024002B303EB025E01D5016E01E4010D02BD0015039602D30206023E00B1025D0389035102F2027B014A01EA021600EA02360143023F01CB0278013402FE014B0367036A03110328032E009301ED014D009F00B7035A0260018D02BC033401580036014401B90133018800BB030E027A00460037022000DA0003018C028F021803B40001017500AD0246014803CA01DE017603E601DB033F03D8024E02CF006302CD001D01FE02C801BE03160338033B024D0298008902770314003C01BD00EC,16384'h003400970025021E038F01AB01F602F602F702410161006202120328027D018802750047001302A100E7000503CF02E000AF021600260213008400A6038B022300C5034702CE0200019000A1028D031C033C021501D4030B0094019E03C00184010101F0004C01990388024E0398015202B800BA028F02C700A5008A03100166036002B9002D03C601A0001603610041001400F70070002E03C2019D03DA01BF02BD020F036301CE03AD0321011E037103BD028C01B500C20367014302B3001D01A1012D015D005802AB007F007803300320034F0024039A0142029F030103E0020500A3025001CF00DA001B031700DC0196012003BC0279011C001E01A6005A02B7017000AE03C702C3034B031D00FD010202B003D800FA03AE0240039401D90057023D023502B5007502E8032B017300E50002025D0195020202EC006F018F010801D6029403DB0137000100E3030803B300E103A801B100B402F403DF0011026400810217018900D90314002B005F0091031502EE01FE0253035B02F10093035703FC012100DE027C022701AC03CD00D701930322014B0124010E010F03D7001000ED0280030401B80267020900B0005E03A000F802710369019201A400E2003503790004039E02D5039C0175014A00CC01E300CA02FD00DF00B7015503C1012B0285033203F8016E015C0286025F03D203650146011001C7034D005B010C03EE03F701630187013902EA038E01600274037B026C00A4009E02B102780287031F007901BD000D006103F0033B03B0025902CA0312001A00630229014F03D6017C011401E2004900B801DE00FC01E7010D00F0017F03C50106038403B503B8039201D7018D030001DA00F6021101C00052025E02B4011D00B3037C02B6009F00BD0219018303ED0126024A0007005D003B008B03B2034A03CA011B01F402DA00CE022E037A016B01F301C403CE0179013D0172016203FF033102490150030A007B03EF014801E1012901BA00EB02E2029602E402470341033D025A006B006001FA009503330045015E038900FB01AE032302EF0036014101B700B2018B0319003703A90343018002AD039702260092023C02D101C8033F022C00F30027036803A601350044019101810178022A019A01DD007401650244014700BB032A01FF03640033027302EB0255019C02C9037F008F03A50383011803DC02D201B302DD00D3016F0238034201E0030702240214029D02F200A00031023A032E03A200F4005300F50116031B034E02D403D3002C03E200BF02820220033A038103AA009A009901B402C1006801FC03EC013C0122010A027B01E6023E02AF0385009801CA0042033400B5036E02B2004A029A0346037500D602A601C1020E007D00AA01D000BE016D026D020403EA014C01850362004301BC019B015F00F9035C01C301000089032D01B20176030F02680348033E00E001A30354035A03900109018A02AA01BB0393024C03050009036F02BF02AE025B03E30376034401C200A2007302610326013A0254039D00290086015701EB0208022B00AC02BB003801AD0269021A035D01B901B6009B026B01250327010700EA014E0000011F03CC00B90339013800A702DE00FE02E503F601F7009C015302D00140004F033800300270000F0131025C03FB0231038A00E6007703B9001903FD002F03E7023601A2039B000803EB00D50096015100CF01ED02BC024B017B01940257021B008200C903D1034C01EA0246037201A80291012700D201A5007201EC03C403DE02CB00AD0353026502A802E3006C03D502D9001203A30111037703FE022800870198003C03CB026303A4005100F102C401EF00E40136029E0182007100DD01D300E903F3029703C300C4009002F900C70266026F037803BE023401F903B700EE02CF036A035002F5006A0021020C039601F102C50352029501BE00690048030D00C601C5014400EC02E103C902E90022006603E901AF03B600A8006402AC000600FF02DB01EE0028023F0391003F003A01F800C80123031E03E4032F01680309001702D3008302320248034500B603FA02F001DC011202D6010B012E029C007C02A3000E02BA0260028A0370019F01E900E803B40222032C005503F100C1001501E402890003005002F3009D0203011A03D9013402D801CC02A2036D028E02A402CC01FD02FB02DC029001D100CB021801E8018C02A9004E021C016903D400B103990018008E027F01D501D8026E02C6029B02430159011901450373037E00D40395038601030374005C02C8017102FC01CD008C0023015800BC020601050177038C036C0258005402FF022D0283016C03820132007603180040031100CD030C02FA002A017E022501CB01A7013F00D002520032037D00D1001F024F02C20284027E026203560221012C023B03370113000C03DD02A0013300C3013B0306003E006D006E016A001C02A70237003900850351033603A101FB03F5021D03AB01B003BF02CD014D0358026A01970272008D0128029203E8005603590230017A020102FE017D0207024201DF032502F8007A00EF01300329030E01C60233014901C903F2013E0276020A02A5015603F9012F03E101D200DB03BB02E703A700A903E6024D020B025600800154011503AF004B00AB03B100C0036B028B018E03AC02C0000B0316027A035E0088033501F200D8007E0324027701DB03C803BA0065011700F202DF0387034903020245015A0313038D006702ED02930281023903400164021002E6031A0366035503F400460288005901AA0299003D00200380010403E50167035F01A90174015B03D0000A0251022F020D012A01E502BE021F0186029802D70303004D01F5039F,16384'h017C026800FA0367007203C00142035900730112037103FD02FE02E6038303110012000F0277022B023D001E032F0291020300CA02AB00D901B8030500CE015601D40094031D01BA01C8011D032D00D6028903C4031503EB00AF0368004501C703F402B100590027033801B5021F030D021C0143027E028601D503730280028103D300E600E202430062026101A7029C0071020E0333018500EC01F703EC02A50107015C03DA0008000D017A00A00129008203D802E201BE03FE00FE025B038E016B01F003E30043035C037D00BD001501030384030302A902D0018E039F0201017402BC030F0312014103B90332030B025202D3022401D0006E008C021400DF006D019C03250250039D03A702AC03C302ED004802DF01DD03C602D801EF00B901930041032101F403BF00D00067023C016101D2020001CE007C00D102E7003F017502C801AC031B000C03C1029D026B038C03C5016603F0003502F203B203E001A20238039102FA0117003000F60320030A023B0381028D027800E9034A03A20202037A001900CC01D60036005B0390015802DC016A001300FF01A902A802D60046010E025E01E8018401380218018A0162013C03DD0331030002870115025C03A4033602B6032E01A003FA004E0011036502AD02D4028E02C901E003CE009A01C5015200C0012302AE002B00A503610272019402FF02CF01A802EB01E60340012E01DC0309034C02F302D702A7039E000101360157023703BE03C9016901800349026C0078036B02E9022000F9009001D300B302DA01BF032201F601FA00BC031000B102EF0344009D025D002E03C802990360028B02BB014803B402E8013B0207013902470050012C01FF02D5032A003901000055027F038703CF0229012401440121024002F001F803D602B70324020A026F0330002C03BD0037038800B70236021200FB007002A20085022A00A1032C01ED027402C30258005A010B025A03DF037B01250295001002F500310347001401500394009600AD012701EE002602BA01BD00AC012F0328004402EA0329021B01EC0262009500D500CD0189007B02930209030701BC020C03E601A103CB01EA018C0060004B019B03AE010A02A4019501770350021003BC005D02630176006503D701A3007D00D2028401AA0251013103F9020803E20267038A0058003400BB0341034603D2007A0128033901180149008002410366033F01B9021A01110259039202F6008D02830171024A011E020400C8014501FD001803EE01FC027C02AA03270282021300DC016D037E002A010D022F011001260215038F009E038D016C00D403F80049011F01AD001D01E203A602310270007F0061039A00BA03AD03450020030801E103A503B7005200B0001C021103EA0079039B02F1003D033A018B00AB005102B000400230013A026D01BB004F017303A103AF0374035E03D103CD015D02DB004C0057021D02EC005403040362009200A900DD0370013F02B9015100C40227022502C6037F006C035400890042010C0159019D0006015B002402A30269006300FD0003016E015503930378010100EA00E50314015E002901DE0033034D03F602E102F901CB02BE03FB020F008701200244008E035A00EE00C3016F01E4013400DB00C601AB028A00F401B302C4000E035D014D01D7027902B5007E006A012D002D032602B403ED000A0098008303C70190024F02DE03DB003E00F801E301D8008B023F03B000CB00D70097015F022D03160228027D00D800B203AC025F0232002202D100F0014C008F0005003C00E3025303A902EE03E5028C0337003B010603E10047029B00280183023E007600BF006401AE0032026E018F00B800C103E703750122027A024B025500D30242001F03820109012B0364016803E400A803BB033B0086014702C5022601EB036901CF001A01CC03AA00E702B80104023303CC0199034301B0008803E9033402C0035800C503EF028F01C601CD02BD011C01A500F1036E031F01A6004D00C2029702210160019A00A200E800E000F20294020D006F036A019201C103B8031E0165013703C2010200A702DD011601B6030E033E02F803D003190009035500B603B501C4039C008A0248012A01FB01CA039503FF037C013E00380352008100A30186014A02E301D902A1019F005602FB03F300DE0385018D0372034E037601E901C0026000EB0007032301B1009B0363009C02340245001B00F7017903DC0256011A009F033D00DA015A005E01C301F1011301910130024E03BA0178002F017B00F500680197023A017F0188020601D1035B0348000202F400170265038B02CE01FE027501A403E801810389030C029A01B700E402A002C7021701F3014F038601B200FC01E503010239013503B30091024C013200E100B501870379032B0276027B02CC021900B4027302CA03990105017E03060093034202C202D2002502BF03B601B40290036D02CB034F03510154017002FD03A3011B000B036C02A602F7033C014002C1010800A6017D0292024D02AF02B3009900BE03CA039703F5021E00530182027102E500210317022C01C9035601F501F2013300CF029F0172014B00AE00C901AF005C01E7004A034B03A000F30296000003D502220119010F0223000403350114029E00ED0216006603AB00AA003A007701DF0198016401DB0249031A0254019E03180153005F0075007403F2014602B2014E022E0257037703FC00C700A40167013D03D9026403D402E00298039802CD03800235006B01DA028502E40069039603020357024603F700EF02FC03DE01F900840023035F03F1031C0016020B03B1026A019601C20205036F0313016302880266035303A802D9,16384'h0020032F0384032B01BE002A011F006201840214039C0085030A031C035600FD01AC03A501140385022D01DD02FB015F02DF0258023201BF011E01D503BD03C70279035A007402C001750317011502C601CF0221023600E0018E012E023F018B0141013703EF015A025600D6037103CB03DD012801B1015D016B036A00BC020C02E801CA029A02EF0055022303C00182013E00ED039400970004018302F10286010003E6024D008703AA01AA03C603C202B9014202E702AD00BD0329022B02FF01C902C8034B028F02BC00020204020E038900B1011803B3029603F2031F0351011301BA0076019000D300FB01500071038301E000EE02920127027C00F001E200D700820310020B02BE02E102B500D501EE008F00B50272004103E403EC021500A7014A021801A6007901C50208022F0084039802A500DC02450045004D004302F900CD037503F80044031803AD016C00CC01040158008C002102F703B000F403570033021E026D0092038002A8004A003E03DE032702CE00E801A9013503BE0255019D02AB004B038E0237007C037D006900420101039D03E80073029F00030302008D00AA03E302250178025C0344036600AE0106010D00C0035D0257032102F2000D005601BC014902AF033D032E021201FA0319032D0283035203C101FD01FE01E503CD0303009E0350025F0275003F03F9029802A3015C03A103F4032800C90370025903D702DB004C005B007A02A00013033E01F9037F03BC00C3027102A6026501DF015902B20388000C03A30289001D016F034F031603DB0179037B010C01BB014600DD0086023D02E0005A029402A2017B00DA00DE004700A802A103AB03D0024800FC02110374000103FA015E034201F0012901E401C1017202FC010E005803B4005F01F1036B0040010A009B01BD009C019600B7017A026F0133019101CD0122001703EE03FF001C002203A602D5036C01470064025D028A0199033500240315010702B00038033F0220028B0132029900BF031D02B7019702B800BE02F802A400A0036400000121037E038C0186031B00F1000A0334013603B800C4033000E3038A03D602AC01DB002B0227005301CE004602DC008B017E02C3033300E9016E0139006A019F01E702E4029501EA028203FD03E0026E00290373009303B7031E00F5022A022C03250381035B018A01EF002C024201FF035C02CB0091023C03AE00A3039E012D00EB01B40034023502EB0205033101F502C703CA025A028700C20168014E01A20189000803FE0217006C0065001102EC019C013002D101F202E202F0021F02880268004E000B0369019A02000311003C001603DF02DE0134013A026100A5015203650009010F00A202440066034103F703D303E9037A00B600940039039601B3038F00BB003201A401C603D1001903D403F3027703E5001E028C001A039001F600B400D2012A01560140020200FE00BA020301B900C5028E011D030E0108021003E2004F03A0034C01A801E900FF026C00A1019E01CC02CA025B033B03DC0154018C03FC03D5019B002603C5033C0006034801B200E5030602C2027A038202F301B601F701ED014400A6016400F9012F036D0397033A02410072013C0143030102F600230320026203ED0353018D01C8038D020A0167005E00EF0054031202E300D1005C0222036F00DB020101D20035037200CA01E1016502460070006E01D0017101AB00CB015103D8003B00F602CC001401E303D2032600D0029E00EC000E014500D902240305019202B30251029C0281023301EB03F6032C0291025201F3036E019801DC014800A4024900E602C901C0017D023903FB0080021C024F024E0018009801FC0273006D03B502C500C802AA033202E601DA03EB00F300B00067023402BF00C603B601D9007F03C400D402FE029303B90307011003CF00B8021A03A203000169034D038701CB016D017F0109029703DA0219008A0355020602160180003D01A100900170009A01A301D400DF02D702DD013D02DA00D8000F026B001B010500F7026603CE014B01B500B201D800B901AF0051004803EA01D70323005D00960181030B024C01C301C20250026000CF01FB018502BA02CD02EE02C1006B0068032A009D0015007801760358027E0247005200E20025012403B100E1039900FA025E01A70103023801730313022900AF002D014C0386009F034E02D402C4005702D602B1028D030C03E102F50037003602A90345021B0125011603B20161031A001F0207016A039A01DE026401D301F400F8015B02D3023000E4034A013100830274024B03D9020902E90077002F020D002E0005026A01230228029B027F016001A003C8029002EA02D80102000702D2013B035E0391011C02D9037C0270015703C30089027603A70267013F027D0155010B029D028000AB02B600C10153034601A50195030F03540361036202400194014F016303BF028401200177002703E7006F039F03360368006002AE003003790187030D034301C401E800120309012B02BD009501B0020F018F016202D000F20263035F0308007D01AE03F10166008E0213012C00590269036000A9014D023102BB02FD01D6019303F503770099027B034901E60081023E01EC0395004903AC03BA022E02ED00EA032202A7036703F003A4011701D101740226023B0028039B007B011B033800AC0363017C0111021D03BB01120188037800B301F8003A024303CC006103C9033903AF013800E7001000CE01AD0314037602E50337035902CF02FA00AD0119006301B8025402F4028503240126011A027803A9008801B7007E0253003100C7034003930392023A030401C70075038B024A005003A8034702B4,16384'h038A03940263016B0052018A036402EC014303450290020103D6026703930254012500AA021F036B01B10238021303E101CC031B013302FF036303B802CE01EF00790141023C0135011B02DA015B01EA01A00322016E03F2003C01F70257022F007E0181005E014B02B902CF013F001701F9024301A1026600C4004A01DB007002BC011401AB003800F401C1022800930080012F00B2019701DA000A03B7000E00BC00C5036F00DD026D023B004D00D0018303BC016F01BC03600205026903E5034200DA03A901370051001901FB023D02D100FC01F5016D03EF017E00090291008403F903EA00ED00C2026C01470219014901A2008203340371032A014D005801D7027503AE029F00A903F4007D02AF000501C902DB039601130091015E014F0248013E031300B40332034C03260014009200F6011801E60016034E01E100FB033302A50308029303300169022201DD02BD01240236039A0325033D01EE0111023A030203F7013803F600FE02B203C002840123039E00C10386017C0086001502A100EF0298024F00B9010902060357033B0060012B0026034302D000C603050397003402390359026E03FA0077039C035D011A037E0288035E028B032B0174013A025A025E02990338028D008B034102FB00D603DA02650249009F00E5018001E200BB020E0235009A014C01AC009703AD033F00E1007B032700A601FC03F3000C028E01C801FA009803360203011C006100B7001302EB0020014E006E038302C5028101B60349003D020400A80395004103EE00540002019000FD039F022303BA0226029400940323024C028C020C01DE002400760362001103CB029E031E006601B9037D01A500AB008803A201E001E3006C000403D400BA00BD0369037901B3012E01CD023001B800B803E7022402FD02C200D2036E002F02C8030900A7027C0139035C021A027E013B02A6015202D7036502CA0384030301F600FF02760157025600D402C401F401750173018D037C03C2006B03FB004B009E02AE03CF03C100CE02B70101025C011F031F020903D500B6024B012001B0018E01CE02D2030B019E036A005F030401CA035600E4016302DE00960108002C02C603A603210031011600CA02EF00E00261022E0368039D0273021200450399001A02F60112006800E6029203BE005302C903B503AC03DF02AC038F03CA025800F000C802B60006027101BA00280355017F03580244034F00DF0354035F039200EA01270240037201A6005A020A015902E0007A019A004701A90110009003B60172013603A7029B039101AD02DD038E027F03E3018201910390010D034A013C015603C7006A03F1031A00AD028201C0037A01AA0010004201C4011503F503F0021B001C023402080280019903A0030702A302E202B103C602F002520231007103C3020D039800740107030003FC01D103DC021403E803A1010E01760278032F012101DF02FC00E801BB0195031C036100670087036D03BD038C027B015F028A008E003E0142038902A703E401BF03E902E7021C02A200D802B30253019B026002F803A8004401A4009B02BE032E0262033A03FE0037035A02E5012601BE029603B400CB021100F303E2027D01A7024602EA006202E300630105037803B903D7033102C1018702C302F202E902F7012A007C0344028F0186010A01CF027003D000640188005B021601B5019803A30388013D03400374038B00A10056020202950145014A0158018F01960075000801E903C8004601610329024502A0009D02510085030F016602F302830128021003E603C5022B01F200F50315002700DB01BD019400EC03EC02000089035302F4022501D9015C01AE0083018902CC0131035103AF00D1001E01F1000B006D016000A20350022C00E903BF0227023E0207036C03A4022A001202E401E403ED00D300C3010F02D902A80153015A00DC004902B80179016501E7003001EC01F80277030E035B030C00CD03D3033903AB03870250012C023F02FE03BB00EE020B031D0221009501B70177004E02AB012902D60104018400E701FD01320312039B01E50148008F037F0242001F034D0306011E007300A4024700070335021803EB027202EE03670348007800D90347024E01920317016800BF02D303AA03DE0033031802E8026B026F024A00F80170025901ED01D400E301C60100034B00F202C00022003F02F500D502790072008D029A001B0171010201B400210154016701AF033C03FF03D101E8035202C7015D0382021D017A0164011D03D8009903010268021E02B5013403E000B1004F02410274006F002A00DE024D01C70039031102DF02AD00F9028700B50264032C03C401DC03B003CE037B0346002B019D02A9009C015001C200A5032403B3023202F900B30144032801D20185004C016C02AA03CC02E100CC005903D2002900FA0297003B03D902B40043025B0314022903F80119004002200023005702D403CD011703660032029C0286037701780215032001B201D5037502D80069012D008A0370025D033E006502CB016A037603B101EB00BE0233010C01A30025008100EB004803A5005D0193005C010B02BA01A8022D00C0018C028500F7038502BB02E6008C0162028903DD027A01FE00E2002E02ED025F017D000F01D003DB019F00AC018B03B2001D01C502CD00AF0001029D007F00CF0310020F01220140019C03C90337002D021703FD01C300C702DC02FA030A01300373003A01D60000026A00A3010601D301FF030D00AE02D501F300A0003501D80255003602BF00B00155038000F1010301CB0319017B015100030237001802B000D701F0038D00C9032D02A4000D0381005500500146031602F1};
  

  genvar i;
    generate
    for (i = 0; i < STATE_SIZE; i = i+1)
    begin : loop1
       assign next[i][0] = {sbox2[i][(in[(i*64+6)+:10])*16 +: 10],sbox1[i*4][(in[(i*64)+:6])*8 +: 6]};
        assign next[i][1] = {sbox2[i][(in[(i*64+22)+:10])*16 +: 10],sbox1[i*4+1][(in[(i*64+16)+:6])*8 +: 6]};
      assign next[i][2] = {sbox2[i][(in[(i*64+38)+:10])*16 +: 10],sbox1[i*4+2][(in[(i*64+32)+:6])*8 +: 6]};
        assign next[i][3] = {sbox2[i][(in[(i*64+54)+:10])*16 +: 10],sbox1[i*4+3][(in[(i*64+48)+:6])*8 +: 6]};
      
      assign out[`IDX64(i)] = {next[i][3],next[i][2],next[i][1],next[i][0]};
    end
  endgenerate
endmodule


module odo_apply_masked_swaps(input [639:0] in, input [639:0] mask, output [639:0] out);
  wire [639:0] swpin;
  assign swpin = {in[`IDX64(8)],in[`IDX64(9)],in[`IDX64(6)],in[`IDX64(7)],in[`IDX64(4)],in[`IDX64(5)],in[`IDX64(2)],in[`IDX64(3)],in[`IDX64(0)],in[`IDX64(1)]};
  assign out = in ^ ((in ^ swpin) & mask);
endmodule

module odo_apply_word_shuffle_rotations(input [639:0] in, input [39:0] rotation, output [639:0] out);
  localparam PBOX_M = 3;
  localparam STATE_SIZE = 10;
  genvar i;
    generate
    for (i = 0; i < STATE_SIZE; i = i+1)
    begin : loop1
      assign out[`IDX64(2*i)] = (in[`IDX64(2*i)] << rotation[`IDX8(i)]) ^  (in[`IDX64(2*i)] >> (8'd64 - rotation[`IDX8(i)]));
        assign out[`IDX64(2*i + 1)] = in[`IDX64(2*i + 1)];
    end
  endgenerate
endmodule


module odo_apply_word_shuffle(input [639:0] in, output [639:0] out);
  localparam PBOX_M = 3;
  localparam STATE_SIZE = 10;
  genvar i;
    generate
    for (i = 0; i < STATE_SIZE; i = i+1)
    begin : loop1
      assign out[`IDX64(PBOX_M * i % STATE_SIZE)] = in[`IDX64(i)];
    end
  endgenerate
endmodule

module odo_apply_pbox_rotations(input [639:0] in, input [39:0] rotation, output [639:0] out);
  localparam STATE_SIZE = 10;
  genvar i;
    generate
    for (i = 0; i < STATE_SIZE / 2; i = i+1)
    begin : loop1
      assign out[`IDX64(2*i)] = (in[`IDX64(2*i)] << rotation[`IDX8(i)]) ^  (in[`IDX64(2*i)] >> (8'd64 - rotation[`IDX8(i)]));
        assign out[`IDX64(2*i + 1)] = in[`IDX64(2*i + 1)];
    end
  endgenerate
endmodule

module odo_apply_pbox(input [639:0] in, input [640 * 6 - 1:0] mask, input [40 * 5 - 1:0] rotation, output [639:0] out);
  localparam PBOX_SUBROUNDS = 6;
  wire [639:0] process[15:0];
  assign process[0] = in;
  genvar i;
    generate
    for (i = 0; i < 5; i = i+1)
    begin : loop1
        odo_apply_masked_swaps swaps(process[i * 3], mask[(640 * i)+:640], process[i * 3 + 1]);
        odo_apply_word_shuffle shuffle(process[i * 3 + 1], process[i * 3 + 2]);
        odo_apply_pbox_rotations rs(process[i * 3 + 2], rotation[(40 * i)+:40], process[i * 3 + 3]);
    end
  endgenerate
  odo_apply_masked_swaps swapst(process[15], mask[(640 * 5)+:640], out);
endmodule


module odo_apply_rotations(input [639:0] in, input [8 * 6 - 1:0] rotation, output [639:0] out);
  wire [639:0] process;
  wire [639:0] next [6:0];
  assign next[0] = {in[63:0],in[639:64]};
  genvar i;
    generate
     for (i = 0; i < 10; i = i+1)
    begin : loop1
       assign next[1][`IDX64(i)] = next[0][`IDX64(i)] ^ (in[`IDX64(i)] << rotation[`IDX8(0)]) ^  (in[`IDX64(i)] >> (64 - rotation[`IDX8(0)]));
        assign next[2][`IDX64(i)] = next[1][`IDX64(i)] ^ (in[`IDX64(i)] << rotation[`IDX8(1)]) ^  (in[`IDX64(i)] >> (64 - rotation[`IDX8(1)]));
        assign next[3][`IDX64(i)] = next[2][`IDX64(i)] ^ (in[`IDX64(i)] << rotation[`IDX8(2)]) ^  (in[`IDX64(i)] >> (64 - rotation[`IDX8(2)]));
        assign next[4][`IDX64(i)] = next[3][`IDX64(i)] ^ (in[`IDX64(i)] << rotation[`IDX8(3)]) ^  (in[`IDX64(i)] >> (64 - rotation[`IDX8(3)]));
        assign next[5][`IDX64(i)] = next[4][`IDX64(i)] ^ (in[`IDX64(i)] << rotation[`IDX8(4)]) ^  (in[`IDX64(i)] >> (64 - rotation[`IDX8(4)]));
        assign next[6][`IDX64(i)] = next[5][`IDX64(i)] ^ (in[`IDX64(i)] << rotation[`IDX8(5)]) ^  (in[`IDX64(i)] >> (64 - rotation[`IDX8(5)]));
     end
  endgenerate
  
  assign out = next[6];
endmodule


module odo_apply_round_key(input [639:0] in, input [15:0] roundKey, output [639:0] out);
  assign out[0] = in[0] ^ roundKey[0];
  assign out[63:1] = in[63:1];
  assign out[64] = in[64] ^ roundKey[1];
  assign out[127:65] = in[127:65];
  assign out[128] = in[128] ^ roundKey[2];
  assign out[191:129] = in[191:129];
  assign out[192] = in[192] ^ roundKey[3];
  assign out[255:193] = in[255:193];
  assign out[256] = in[256] ^ roundKey[4];
  assign out[319:257] = in[319:257];
  assign out[320] = in[320] ^ roundKey[5];
  assign out[383:321] = in[383:321];
  assign out[384] = in[384] ^ roundKey[6];
  assign out[447:385] = in[447:385];
  assign out[448] = in[448] ^ roundKey[7];
  assign out[511:449] = in[511:449];
  assign out[512] = in[512] ^ roundKey[8];
  assign out[575:513] = in[575:513];
  assign out[576] = in[576] ^ roundKey[9];
  assign out[639:577] = in[639:577];
endmodule


module odo_encrypt(input clk, input read, input [639:0] in, output reg write, output reg [639:0] out);
  
  wire [640 * 6 - 1:0] mask1 = 3840'h66E8107925D7FE0966E8107925D7FE09C25CD32259AE83CEC25CD32259AE83CEFD23D04576C7734EFD23D04576C7734EA34AADDF49D8DE64A34AADDF49D8DE647D91DEB549A4F1477D91DEB549A4F14715F5C877017BC76E15F5C877017BC76E9B7F04D1BAF2C4699B7F04D1BAF2C4693FFE91D3446F4C5C3FFE91D3446F4C5C6436019CE44360676436019CE4436067440EDCD2076DEA01440EDCD2076DEA01D74B878A9643DDBFD74B878A9643DDBF25A4BF2D4B3D2C3D25A4BF2D4B3D2C3D72EE006070AEBA7D72EE006070AEBA7DAD4A08AFF581F5B8AD4A08AFF581F5B8DBA44032C2BF27D4DBA44032C2BF27D454D60DE2E96CE37854D60DE2E96CE3789CC4EE726ACC72559CC4EE726ACC7255AC060DC1CA4BB5C6AC060DC1CA4BB5C6843A1E2F68208610843A1E2F682086104CF5A158B7B702604CF5A158B7B70260217B3CCF03E49E73217B3CCF03E49E73F7A1062DD1C651B6F7A1062DD1C651B686E11CD92075461186E11CD920754611BC68536E2A668DDDBC68536E2A668DDD67FC1EBCA60F57B267FC1EBCA60F57B2F1474338BC7DBC92F1474338BC7DBC9232169F07D2028A4932169F07D2028A49887855B94F175C50887855B94F175C50C566AC13A7D3DADEC566AC13A7D3DADE74392302F726B2DC74392302F726B2DC;
  wire [40 * 5 - 1:0] rotation1 = 200'h2D1811093B0C2A11292B1A323A1808080F26011D3C0F3D3708;
  wire [640 * 6 - 1:0] mask2 = 3840'h48801E29D10E7B8048801E29D10E7B8002674114B6AEDE4002674114B6AEDE40EAECA60D4502A639EAECA60D4502A639D7AA3DF885A8D3BBD7AA3DF885A8D3BB03CD28179848F24D03CD28179848F24D8B5B954A69FFA9618B5B954A69FFA96151A8BC89F40F6BDD51A8BC89F40F6BDD426F7EC429FA4D41426F7EC429FA4D4186A5AD69C7496A0986A5AD69C7496A09B4050C921732716BB4050C921732716BDC4C64FEC218343EDC4C64FEC218343EE010AF61F44F59F7E010AF61F44F59F7F48E75366674C18BF48E75366674C18B4BEA2540C051CDB34BEA2540C051CDB3C9F67094A1777AC5C9F67094A1777AC5F5BFB82DE1046F00F5BFB82DE1046F00A9A625464D32134CA9A625464D32134C0B3B90772827A7EF0B3B90772827A7EF943E5A20BD22183B943E5A20BD22183B7A86D20B31B1C5867A86D20B31B1C5863DE8D7F3D09D948C3DE8D7F3D09D948C4B079C4EE95969334B079C4EE95969339B996D2562B013729B996D2562B01372E0DD9520A929733BE0DD9520A929733B6793F75AB3B754216793F75AB3B754216B8D8C52D70D44556B8D8C52D70D445537E76087C49C094837E76087C49C0948758DB972CA844A19758DB972CA844A194F45686CF2D2A5204F45686CF2D2A520526CC04FBCC86390526CC04FBCC86390;
  wire [40 * 5 - 1:0] rotation2 = 200'h2E0B3505361F1A031C27140B2E13293322393614311E101D0B;
  
  wire [8 * 6 - 1:0] rotation = 48'h052709371732;
  wire [16 * 84 - 1:0] roundKeys = 1344'h01FD01DD03DF02F0020402C300C80104026702050132032903F3016503F000E90148032D008403F7028C00060188017C031F004F0000014F0286025E0087039E0102035002E6008E03F70024008401850048036502B400EA01B500BD02520226025901FF039302DF010603E3036D017E03E900DB02C0039601D2010502F20026010901C900170167021B02EE039B003B01C9000B012402E900AB01CF030A00C90051001F013201A3;

  
  localparam ROUNDS = 84;
  wire [639:0] process [5:0];
  reg [639:0] data;
  wire [639:0] mixdata;
  reg [7:0] round;
  reg[15:0] roundKey;
  
  assign process[0] = data;
  
  odo_pre_mix mix(in, mixdata);
  odo_apply_pbox pbox(process[0], mask1, rotation1, process[1]);
  odo_apply_sboxes sbox(process[1], process[2]);
  odo_apply_pbox pbox2(process[2], mask2, rotation2, process[3]);
  odo_apply_rotations rotp(process[3], rotation, process[4]);
  odo_apply_round_key rk(process[4], roundKey, process[5]);
  

  // 开始计算
  reg [1:0] cpstate;
  always @(posedge clk) begin
    cpstate <= {cpstate[0], read};
  end
  
  always @(posedge clk) begin
    if (cpstate == 2'b01) begin
        data <= mixdata;
        round <= 8'b0;
        write <= 1'b0;
        roundKey <= roundKeys[15:0];
     end
     else if(round < ROUNDS-1) begin
       roundKey <= roundKeys[(16*(round+1))+:16];
        round <= round + 8'b1;
        data <= process[5];
     end
     else if(round == ROUNDS-1) begin
       write <= 1'b1;
       out <= process[5];
     end
  end
  
endmodule